library verilog;
use verilog.vl_types.all;
entity tb_vga_ctrl is
end tb_vga_ctrl;
